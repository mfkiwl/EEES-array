////////////////////////////////////////////////////////////////////////////////
//                                                                            //
//    Module Name :  simd_top_testbench                                       //
//    Description :  Template for the testbench for the SIMD processor.       //
//                                                                            //
//    Author(s)   :  Yifan He                                                 //
//                   Dongrui She                                              //
//                                                                            //
////////////////////////////////////////////////////////////////////////////////

`include "def-cp.v"
`include "def-pe.v"

`include "def-testbench.v"

// synopsys translate_off
`timescale 1ns / 1ps
// synopsys translate_on

module simd_top_testbench;

//******************************
//  Local Wire/Reg Declaration
//******************************

  reg                                   rClk;   // system clock, p-edge trigger
  reg                                   rReset; // global sync-reset, cctive low

  wire [(`DEF_CP_I_MEM_ADDR_WIDTH-3):0] wPC;      // PC to indicate the end of the program
  reg  [(`DEF_CP_I_MEM_ADDR_WIDTH-3):0] rLast_PC; // buffered last PC
  wire                                  wTask_Finished; // self-jump, indicate the end of the program

  // instruction memory
  reg  [31:0]                           CP_IMEM_Init[0:(`DEF_CP_IMEM_SIZE-1)];
  reg  [31:0]                           PE_IMEM_Init[0:(`DEF_PE_IMEM_SIZE-1)];

  reg                                   rBus_IMEM_Valid;       // ins. memory access valid
  reg  [(`DEF_CP_I_MEM_ADDR_WIDTH-3):0] rBus_IMEM_Address;     // ins. memory access address
  reg  [(`DEF_CP_I_MEM_ADDR_WIDTH-3):0] rBus_IMEM_Address_Next;// NEXT ins. memory access address
  reg  [63:0]                           rBus_IMEM_Write_Data;  // ins. memory write data
  reg                                   rBus_IMEM_Write_Enable;// ins. memory write enable

  wire [(`DEF_CP_INS_WIDTH+3):0]        wBus_CP_IMEM_Read_Data;// cp ins. memory read data
  wire [(`DEF_PE_INS_WIDTH+4):0]        wBus_PE_IMEM_Read_Data;// pe ins. memory read data


  // data memory
  // CP
  reg  [(`DEF_CP_DATA_WIDTH-1):0]       CP_DMEM_Init[0:(`DEF_CP_DMEM_SIZE-1)];       // CP data memory
  reg  [(`DEF_CP_DATA_WIDTH-1):0]       CP_DMEM_tmp[0:(`DEF_CP_DMEM_SIZE-1)];        // tempory buffer for dumping cp memory data
  reg  [(`DEF_CP_DATA_WIDTH-1):0]       rCP_DMEM_Reference[0:(`DEF_CP_DMEM_SIZE-1)]; // CP reference data memory (for debug only)

  reg                                   rBus_CP_DMEM_Valid;                       // cp data memory access valid
  reg  [(`DEF_CP_D_MEM_ADDR_WIDTH-3):0] rBus_CP_DMEM_Address;                     // cp data memory access address
  reg  [(`DEF_CP_D_MEM_ADDR_WIDTH-3):0] rBus_CP_DMEM_Address_Next;                // NEXT data memory access address
  reg  [(`DEF_CP_DATA_WIDTH-1):0]       rBus_CP_DMEM_Write_Data;                  // cp data memory write data
  reg                                   rBus_CP_DMEM_Write_Enable;                // cp data memory write enable
  wire [(`DEF_CP_DATA_WIDTH-1):0]       wBus_CP_DMEM_Read_Data;                   // cp data memory read data

  // PE
  reg  [(`DEF_PE_DATA_WIDTH-1):0]       PE_DMEM_Init[0:(`DEF_PE_DMEM_SIZE*`DEF_PE_NUM-1)]; // PE data memory init
  reg  [(`DEF_PE_DATA_WIDTH-1):0]       PE_DMEM_tmp[0:(`DEF_PE_DMEM_SIZE-1)];     // tempory buffer for dumping cp memory data

  reg                                   rBus_PE_DMEM_Valid;                      // pe data memory access valid
  reg  [(`DEF_PE_D_MEM_ADDR_WIDTH-3):0] rBus_PE_DMEM_Address;                    // pe data memory access address
  reg  [(`DEF_PE_D_MEM_ADDR_WIDTH-3):0] rBus_PE_DMEM_Address_Next;               // NEXT data memory access address
  reg  [(`DEF_PE_DATA_WIDTH*`DEF_PE_NUM-1):0] rBus_PE_DMEM_Write_Data;           // pe data memory write data
  reg                                   rBus_PE_DMEM_Write_Enable;               // pe data memory write enable
  wire [(`DEF_PE_DATA_WIDTH*`DEF_PE_NUM-1):0] wBus_PE_DMEM_Read_Data;            // pe data memory read data

  // control signals
  reg                                   rProgram_Finish;                // is the last instruction

  reg [31:0]                            rTest_Counter;                  // data counter for debug
  reg [2:0]                             rPlace_Holder;

  wire                                  wCore_Reset;                    // core reset signal

  reg                                   rIMEM_Configure_Done;           // IMEM initialization done
  reg                                   rCP_DMEM_Configure_Done;        // CP DMEM initialization done
  reg                                   rPE_DMEM_Configure_Done;        // PE DMEM initialization done

  integer                               i;


//******************************
//  Behavioral Description
//******************************
  // ========
  //  clock
  // ========
  always #(`CYCLE_TIME/2.0) rClk = ~rClk;


  // =====================
  //  instruction memory
  // =====================
  // configure imem (cp + pe)
  always @ ( posedge rClk )
    if ( rReset == 1'b0 )
      rIMEM_Configure_Done <= 1'b0;
    else if ( rBus_IMEM_Address == (`DEF_CP_IMEM_SIZE - 2) )
      rIMEM_Configure_Done <= 1'b1;
  // end of always

  always @ ( posedge rClk )
    if ( rReset == 1'b0 ) begin
      rBus_IMEM_Valid        <= 'b0;
      rBus_IMEM_Address      <= 'b0;
      rBus_IMEM_Address_Next <= 'b0;
      rBus_IMEM_Write_Data   <= 'b0;
      rBus_IMEM_Write_Enable <= 'b0;
    end
    else if ( rIMEM_Configure_Done == 1'b0 ) begin   // not configured yet
      rBus_IMEM_Valid        <= 'b1;
      rBus_IMEM_Address_Next <= rBus_IMEM_Address_Next + 'b1;
      rBus_IMEM_Address      <= rBus_IMEM_Address_Next;
      rBus_IMEM_Write_Data   <= {PE_IMEM_Init[rBus_IMEM_Address_Next], CP_IMEM_Init[rBus_IMEM_Address_Next]};
      rBus_IMEM_Write_Enable <= 'b1;
    end
    else begin
      rBus_IMEM_Valid        <= 'b0;
    end
  // end of always


  // ================
  //  CP data memory
  // ================
  always @ ( posedge rClk )
    if ( rReset == 1'b0 )
      rCP_DMEM_Configure_Done <= 1'b0;
    else if ( rBus_CP_DMEM_Address == (`DEF_CP_DMEM_SIZE - 2) )
      rCP_DMEM_Configure_Done <= 1'b1;
  // end of always


  always @ ( posedge rClk )
    if ( rReset == 1'b0 ) begin
      rBus_CP_DMEM_Valid        <= 'b0;
      rBus_CP_DMEM_Address      <= 'b0;
      rBus_CP_DMEM_Address_Next <= 'b0;
      rBus_CP_DMEM_Write_Data   <= 'b0;
      rBus_CP_DMEM_Write_Enable <= 'b0;
    end
    else if ( rCP_DMEM_Configure_Done == 1'b0 ) begin   // not configured yet, configure the data memory
      rBus_CP_DMEM_Valid        <= 'b1;
      rBus_CP_DMEM_Address_Next <= rBus_CP_DMEM_Address_Next + 'b1;
      rBus_CP_DMEM_Address      <= rBus_CP_DMEM_Address_Next;
      rBus_CP_DMEM_Write_Data   <= CP_DMEM_Init[rBus_CP_DMEM_Address_Next];
      rBus_CP_DMEM_Write_Enable <= 'b1;
    end
    else begin
      rBus_CP_DMEM_Valid        <= 'b0;
      rBus_CP_DMEM_Address      <= 'b0;
      rBus_CP_DMEM_Address_Next <= 'b0;
      rBus_CP_DMEM_Write_Data   <= 'b0;
      rBus_CP_DMEM_Write_Enable <= 'b0;
    end
  // end of always



  // ================
  //  PE data memory
  // ================
  always @ ( posedge rClk )
    if ( rReset == 1'b0 ) begin
      rPE_DMEM_Configure_Done <= 1'b0;
    end
    else if ( rBus_PE_DMEM_Address == (`DEF_PE_DMEM_SIZE - 2) ) begin
      rPE_DMEM_Configure_Done <= 1'b1;
    end
  // end of always

  always @ ( posedge rClk )
    if ( rReset == 1'b0 ) begin
      rBus_PE_DMEM_Valid        <= 'b0;
      rBus_PE_DMEM_Address      <= 'b0;
      rBus_PE_DMEM_Address_Next <= 'b0;
      rBus_PE_DMEM_Write_Data   <= 'b0;
      rBus_PE_DMEM_Write_Enable <= 'b0;
    end
    else if ( rPE_DMEM_Configure_Done == 1'b0 ) begin   // not configured yet, configure the data memory
      rBus_PE_DMEM_Valid        <= 'b1;
      rBus_PE_DMEM_Address_Next <= rBus_PE_DMEM_Address_Next + 'b1;
      rBus_PE_DMEM_Address      <= rBus_PE_DMEM_Address_Next;
      //for( i = 0; i < `DEF_PE_NUM; i = i+1 ) begin
      //  rBus_PE_DMEM_Write_Data[(`DEF_PE_DATA_WIDTH*i-1):`DEF_PE_DATA_WIDTH*i] <= PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+i];
      //end
      rBus_PE_DMEM_Write_Data <= {
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+127],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+126],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+125],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+124],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+123],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+122],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+121],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+120],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+119],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+118],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+117],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+116],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+115],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+114],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+113],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+112],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+111],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+110],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+109],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+108],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+107],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+106],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+105],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+104],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+103],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+102],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+101],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+100],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+99],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+98],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+97],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+96],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+95],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+94],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+93],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+92],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+91],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+90],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+89],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+88],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+87],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+86],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+85],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+84],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+83],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+82],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+81],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+80],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+79],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+78],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+77],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+76],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+75],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+74],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+73],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+72],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+71],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+70],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+69],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+68],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+67],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+66],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+65],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+64],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+63],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+62],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+61],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+60],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+59],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+58],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+57],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+56],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+55],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+54],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+53],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+52],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+51],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+50],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+49],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+48],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+47],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+46],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+45],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+44],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+43],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+42],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+41],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+40],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+39],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+38],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+37],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+36],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+35],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+34],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+33],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+32],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+31],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+30],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+29],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+28],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+27],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+26],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+25],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+24],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+23],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+22],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+21],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+20],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+19],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+18],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+17],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+16],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+15],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+14],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+13],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+12],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+11],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+10],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+9],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+8],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+7],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+6],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+5],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+4],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+3],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+2],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+1],
        PE_DMEM_Init[rBus_PE_DMEM_Address_Next*`DEF_PE_NUM+0]
      };
      rBus_PE_DMEM_Write_Enable <= 'b1;
    end
    else begin
      rBus_PE_DMEM_Valid        <= 'b0;
      rBus_PE_DMEM_Address      <= 'b0;
      rBus_PE_DMEM_Address_Next <= 'b0;
      rBus_PE_DMEM_Write_Data   <= 'b0;
      rBus_PE_DMEM_Write_Enable <= 'b0;
    end
  // end of always


  // =====================
  // Last Ins. Detection
  // =====================
  always @ ( posedge rClk )
    if ( rReset == 1'b0 )
      rProgram_Finish <= 1'b0;
    else if ( wPC == (rLast_PC - 1) ) // finsh when jump to itself
      rProgram_Finish <= 1'b1;
  // end of always


  always @ ( posedge rClk )
    if ( rReset == 1'b0 )
      rLast_PC <= 'hAAAA;
    else begin
      rLast_PC <= wPC;
      if (wPC == 'h1)
        $stop;
    end
  // end of always



  // ===========
  //   Initial
  // ===========
   initial
     begin
       rClk = 0;
       rReset = 1;
       rTest_Counter = 0;
       rPlace_Holder = 0;

       // read memory initialization files
       $readmemh("cp.imem_init", CP_IMEM_Init);
       $readmemh("pe.imem_init", PE_IMEM_Init);
       $readmemh("cp.dmem_init", CP_DMEM_Init);
       $readmemh("pe.dmem_init", PE_DMEM_Init);

       #(`CYCLE_TIME * 10) rReset = 0; // 10 cycles;
       #(`CYCLE_TIME * 20) rReset = 1; // 20 cycles
       // test the interrupt signal
       while ( rProgram_Finish == 1'b0)
         @ ( posedge rClk );

       #(`CYCLE_TIME * 2)   // 2 cycles

       // dump cp data-memory
       for (i=0; i<`DEF_CP_DMEM_SIZE; i=i+1) begin
        CP_DMEM_tmp[i] = {inst_simd_top.inst_cp_dmem.dmem3[i], inst_simd_top.inst_cp_dmem.dmem2[i], inst_simd_top.inst_cp_dmem.dmem1[i], inst_simd_top.inst_cp_dmem.dmem0[i]
        };
       end

       $writememh("cp.dmem.dump", CP_DMEM_tmp);

       // dump pe data-memory
       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe0_dmem.dmem3[i], inst_simd_top.inst_pe0_dmem.dmem2[i], inst_simd_top.inst_pe0_dmem.dmem1[i], inst_simd_top.inst_pe0_dmem.dmem0[i]
        };
       end

       $writememh("pe0.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe1_dmem.dmem3[i], inst_simd_top.inst_pe1_dmem.dmem2[i], inst_simd_top.inst_pe1_dmem.dmem1[i], inst_simd_top.inst_pe1_dmem.dmem0[i]
        };
       end

       $writememh("pe1.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe2_dmem.dmem3[i], inst_simd_top.inst_pe2_dmem.dmem2[i], inst_simd_top.inst_pe2_dmem.dmem1[i], inst_simd_top.inst_pe2_dmem.dmem0[i]
        };
       end

       $writememh("pe2.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe3_dmem.dmem3[i], inst_simd_top.inst_pe3_dmem.dmem2[i], inst_simd_top.inst_pe3_dmem.dmem1[i], inst_simd_top.inst_pe3_dmem.dmem0[i]
        };
       end

       $writememh("pe3.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe4_dmem.dmem3[i], inst_simd_top.inst_pe4_dmem.dmem2[i], inst_simd_top.inst_pe4_dmem.dmem1[i], inst_simd_top.inst_pe4_dmem.dmem0[i]
        };
       end

       $writememh("pe4.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe5_dmem.dmem3[i], inst_simd_top.inst_pe5_dmem.dmem2[i], inst_simd_top.inst_pe5_dmem.dmem1[i], inst_simd_top.inst_pe5_dmem.dmem0[i]
        };
       end

       $writememh("pe5.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe6_dmem.dmem3[i], inst_simd_top.inst_pe6_dmem.dmem2[i], inst_simd_top.inst_pe6_dmem.dmem1[i], inst_simd_top.inst_pe6_dmem.dmem0[i]
        };
       end

       $writememh("pe6.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe7_dmem.dmem3[i], inst_simd_top.inst_pe7_dmem.dmem2[i], inst_simd_top.inst_pe7_dmem.dmem1[i], inst_simd_top.inst_pe7_dmem.dmem0[i]
        };
       end

       $writememh("pe7.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe8_dmem.dmem3[i], inst_simd_top.inst_pe8_dmem.dmem2[i], inst_simd_top.inst_pe8_dmem.dmem1[i], inst_simd_top.inst_pe8_dmem.dmem0[i]
        };
       end

       $writememh("pe8.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe9_dmem.dmem3[i], inst_simd_top.inst_pe9_dmem.dmem2[i], inst_simd_top.inst_pe9_dmem.dmem1[i], inst_simd_top.inst_pe9_dmem.dmem0[i]
        };
       end

       $writememh("pe9.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe10_dmem.dmem3[i], inst_simd_top.inst_pe10_dmem.dmem2[i], inst_simd_top.inst_pe10_dmem.dmem1[i], inst_simd_top.inst_pe10_dmem.dmem0[i]
        };
       end

       $writememh("pe10.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe11_dmem.dmem3[i], inst_simd_top.inst_pe11_dmem.dmem2[i], inst_simd_top.inst_pe11_dmem.dmem1[i], inst_simd_top.inst_pe11_dmem.dmem0[i]
        };
       end

       $writememh("pe11.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe12_dmem.dmem3[i], inst_simd_top.inst_pe12_dmem.dmem2[i], inst_simd_top.inst_pe12_dmem.dmem1[i], inst_simd_top.inst_pe12_dmem.dmem0[i]
        };
       end

       $writememh("pe12.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe13_dmem.dmem3[i], inst_simd_top.inst_pe13_dmem.dmem2[i], inst_simd_top.inst_pe13_dmem.dmem1[i], inst_simd_top.inst_pe13_dmem.dmem0[i]
        };
       end

       $writememh("pe13.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe14_dmem.dmem3[i], inst_simd_top.inst_pe14_dmem.dmem2[i], inst_simd_top.inst_pe14_dmem.dmem1[i], inst_simd_top.inst_pe14_dmem.dmem0[i]
        };
       end

       $writememh("pe14.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe15_dmem.dmem3[i], inst_simd_top.inst_pe15_dmem.dmem2[i], inst_simd_top.inst_pe15_dmem.dmem1[i], inst_simd_top.inst_pe15_dmem.dmem0[i]
        };
       end

       $writememh("pe15.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe16_dmem.dmem3[i], inst_simd_top.inst_pe16_dmem.dmem2[i], inst_simd_top.inst_pe16_dmem.dmem1[i], inst_simd_top.inst_pe16_dmem.dmem0[i]
        };
       end

       $writememh("pe16.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe17_dmem.dmem3[i], inst_simd_top.inst_pe17_dmem.dmem2[i], inst_simd_top.inst_pe17_dmem.dmem1[i], inst_simd_top.inst_pe17_dmem.dmem0[i]
        };
       end

       $writememh("pe17.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe18_dmem.dmem3[i], inst_simd_top.inst_pe18_dmem.dmem2[i], inst_simd_top.inst_pe18_dmem.dmem1[i], inst_simd_top.inst_pe18_dmem.dmem0[i]
        };
       end

       $writememh("pe18.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe19_dmem.dmem3[i], inst_simd_top.inst_pe19_dmem.dmem2[i], inst_simd_top.inst_pe19_dmem.dmem1[i], inst_simd_top.inst_pe19_dmem.dmem0[i]
        };
       end

       $writememh("pe19.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe20_dmem.dmem3[i], inst_simd_top.inst_pe20_dmem.dmem2[i], inst_simd_top.inst_pe20_dmem.dmem1[i], inst_simd_top.inst_pe20_dmem.dmem0[i]
        };
       end

       $writememh("pe20.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe21_dmem.dmem3[i], inst_simd_top.inst_pe21_dmem.dmem2[i], inst_simd_top.inst_pe21_dmem.dmem1[i], inst_simd_top.inst_pe21_dmem.dmem0[i]
        };
       end

       $writememh("pe21.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe22_dmem.dmem3[i], inst_simd_top.inst_pe22_dmem.dmem2[i], inst_simd_top.inst_pe22_dmem.dmem1[i], inst_simd_top.inst_pe22_dmem.dmem0[i]
        };
       end

       $writememh("pe22.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe23_dmem.dmem3[i], inst_simd_top.inst_pe23_dmem.dmem2[i], inst_simd_top.inst_pe23_dmem.dmem1[i], inst_simd_top.inst_pe23_dmem.dmem0[i]
        };
       end

       $writememh("pe23.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe24_dmem.dmem3[i], inst_simd_top.inst_pe24_dmem.dmem2[i], inst_simd_top.inst_pe24_dmem.dmem1[i], inst_simd_top.inst_pe24_dmem.dmem0[i]
        };
       end

       $writememh("pe24.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe25_dmem.dmem3[i], inst_simd_top.inst_pe25_dmem.dmem2[i], inst_simd_top.inst_pe25_dmem.dmem1[i], inst_simd_top.inst_pe25_dmem.dmem0[i]
        };
       end

       $writememh("pe25.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe26_dmem.dmem3[i], inst_simd_top.inst_pe26_dmem.dmem2[i], inst_simd_top.inst_pe26_dmem.dmem1[i], inst_simd_top.inst_pe26_dmem.dmem0[i]
        };
       end

       $writememh("pe26.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe27_dmem.dmem3[i], inst_simd_top.inst_pe27_dmem.dmem2[i], inst_simd_top.inst_pe27_dmem.dmem1[i], inst_simd_top.inst_pe27_dmem.dmem0[i]
        };
       end

       $writememh("pe27.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe28_dmem.dmem3[i], inst_simd_top.inst_pe28_dmem.dmem2[i], inst_simd_top.inst_pe28_dmem.dmem1[i], inst_simd_top.inst_pe28_dmem.dmem0[i]
        };
       end

       $writememh("pe28.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe29_dmem.dmem3[i], inst_simd_top.inst_pe29_dmem.dmem2[i], inst_simd_top.inst_pe29_dmem.dmem1[i], inst_simd_top.inst_pe29_dmem.dmem0[i]
        };
       end

       $writememh("pe29.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe30_dmem.dmem3[i], inst_simd_top.inst_pe30_dmem.dmem2[i], inst_simd_top.inst_pe30_dmem.dmem1[i], inst_simd_top.inst_pe30_dmem.dmem0[i]
        };
       end

       $writememh("pe30.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe31_dmem.dmem3[i], inst_simd_top.inst_pe31_dmem.dmem2[i], inst_simd_top.inst_pe31_dmem.dmem1[i], inst_simd_top.inst_pe31_dmem.dmem0[i]
        };
       end

       $writememh("pe31.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe32_dmem.dmem3[i], inst_simd_top.inst_pe32_dmem.dmem2[i], inst_simd_top.inst_pe32_dmem.dmem1[i], inst_simd_top.inst_pe32_dmem.dmem0[i]
        };
       end

       $writememh("pe32.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe33_dmem.dmem3[i], inst_simd_top.inst_pe33_dmem.dmem2[i], inst_simd_top.inst_pe33_dmem.dmem1[i], inst_simd_top.inst_pe33_dmem.dmem0[i]
        };
       end

       $writememh("pe33.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe34_dmem.dmem3[i], inst_simd_top.inst_pe34_dmem.dmem2[i], inst_simd_top.inst_pe34_dmem.dmem1[i], inst_simd_top.inst_pe34_dmem.dmem0[i]
        };
       end

       $writememh("pe34.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe35_dmem.dmem3[i], inst_simd_top.inst_pe35_dmem.dmem2[i], inst_simd_top.inst_pe35_dmem.dmem1[i], inst_simd_top.inst_pe35_dmem.dmem0[i]
        };
       end

       $writememh("pe35.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe36_dmem.dmem3[i], inst_simd_top.inst_pe36_dmem.dmem2[i], inst_simd_top.inst_pe36_dmem.dmem1[i], inst_simd_top.inst_pe36_dmem.dmem0[i]
        };
       end

       $writememh("pe36.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe37_dmem.dmem3[i], inst_simd_top.inst_pe37_dmem.dmem2[i], inst_simd_top.inst_pe37_dmem.dmem1[i], inst_simd_top.inst_pe37_dmem.dmem0[i]
        };
       end

       $writememh("pe37.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe38_dmem.dmem3[i], inst_simd_top.inst_pe38_dmem.dmem2[i], inst_simd_top.inst_pe38_dmem.dmem1[i], inst_simd_top.inst_pe38_dmem.dmem0[i]
        };
       end

       $writememh("pe38.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe39_dmem.dmem3[i], inst_simd_top.inst_pe39_dmem.dmem2[i], inst_simd_top.inst_pe39_dmem.dmem1[i], inst_simd_top.inst_pe39_dmem.dmem0[i]
        };
       end

       $writememh("pe39.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe40_dmem.dmem3[i], inst_simd_top.inst_pe40_dmem.dmem2[i], inst_simd_top.inst_pe40_dmem.dmem1[i], inst_simd_top.inst_pe40_dmem.dmem0[i]
        };
       end

       $writememh("pe40.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe41_dmem.dmem3[i], inst_simd_top.inst_pe41_dmem.dmem2[i], inst_simd_top.inst_pe41_dmem.dmem1[i], inst_simd_top.inst_pe41_dmem.dmem0[i]
        };
       end

       $writememh("pe41.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe42_dmem.dmem3[i], inst_simd_top.inst_pe42_dmem.dmem2[i], inst_simd_top.inst_pe42_dmem.dmem1[i], inst_simd_top.inst_pe42_dmem.dmem0[i]
        };
       end

       $writememh("pe42.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe43_dmem.dmem3[i], inst_simd_top.inst_pe43_dmem.dmem2[i], inst_simd_top.inst_pe43_dmem.dmem1[i], inst_simd_top.inst_pe43_dmem.dmem0[i]
        };
       end

       $writememh("pe43.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe44_dmem.dmem3[i], inst_simd_top.inst_pe44_dmem.dmem2[i], inst_simd_top.inst_pe44_dmem.dmem1[i], inst_simd_top.inst_pe44_dmem.dmem0[i]
        };
       end

       $writememh("pe44.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe45_dmem.dmem3[i], inst_simd_top.inst_pe45_dmem.dmem2[i], inst_simd_top.inst_pe45_dmem.dmem1[i], inst_simd_top.inst_pe45_dmem.dmem0[i]
        };
       end

       $writememh("pe45.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe46_dmem.dmem3[i], inst_simd_top.inst_pe46_dmem.dmem2[i], inst_simd_top.inst_pe46_dmem.dmem1[i], inst_simd_top.inst_pe46_dmem.dmem0[i]
        };
       end

       $writememh("pe46.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe47_dmem.dmem3[i], inst_simd_top.inst_pe47_dmem.dmem2[i], inst_simd_top.inst_pe47_dmem.dmem1[i], inst_simd_top.inst_pe47_dmem.dmem0[i]
        };
       end

       $writememh("pe47.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe48_dmem.dmem3[i], inst_simd_top.inst_pe48_dmem.dmem2[i], inst_simd_top.inst_pe48_dmem.dmem1[i], inst_simd_top.inst_pe48_dmem.dmem0[i]
        };
       end

       $writememh("pe48.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe49_dmem.dmem3[i], inst_simd_top.inst_pe49_dmem.dmem2[i], inst_simd_top.inst_pe49_dmem.dmem1[i], inst_simd_top.inst_pe49_dmem.dmem0[i]
        };
       end

       $writememh("pe49.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe50_dmem.dmem3[i], inst_simd_top.inst_pe50_dmem.dmem2[i], inst_simd_top.inst_pe50_dmem.dmem1[i], inst_simd_top.inst_pe50_dmem.dmem0[i]
        };
       end

       $writememh("pe50.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe51_dmem.dmem3[i], inst_simd_top.inst_pe51_dmem.dmem2[i], inst_simd_top.inst_pe51_dmem.dmem1[i], inst_simd_top.inst_pe51_dmem.dmem0[i]
        };
       end

       $writememh("pe51.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe52_dmem.dmem3[i], inst_simd_top.inst_pe52_dmem.dmem2[i], inst_simd_top.inst_pe52_dmem.dmem1[i], inst_simd_top.inst_pe52_dmem.dmem0[i]
        };
       end

       $writememh("pe52.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe53_dmem.dmem3[i], inst_simd_top.inst_pe53_dmem.dmem2[i], inst_simd_top.inst_pe53_dmem.dmem1[i], inst_simd_top.inst_pe53_dmem.dmem0[i]
        };
       end

       $writememh("pe53.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe54_dmem.dmem3[i], inst_simd_top.inst_pe54_dmem.dmem2[i], inst_simd_top.inst_pe54_dmem.dmem1[i], inst_simd_top.inst_pe54_dmem.dmem0[i]
        };
       end

       $writememh("pe54.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe55_dmem.dmem3[i], inst_simd_top.inst_pe55_dmem.dmem2[i], inst_simd_top.inst_pe55_dmem.dmem1[i], inst_simd_top.inst_pe55_dmem.dmem0[i]
        };
       end

       $writememh("pe55.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe56_dmem.dmem3[i], inst_simd_top.inst_pe56_dmem.dmem2[i], inst_simd_top.inst_pe56_dmem.dmem1[i], inst_simd_top.inst_pe56_dmem.dmem0[i]
        };
       end

       $writememh("pe56.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe57_dmem.dmem3[i], inst_simd_top.inst_pe57_dmem.dmem2[i], inst_simd_top.inst_pe57_dmem.dmem1[i], inst_simd_top.inst_pe57_dmem.dmem0[i]
        };
       end

       $writememh("pe57.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe58_dmem.dmem3[i], inst_simd_top.inst_pe58_dmem.dmem2[i], inst_simd_top.inst_pe58_dmem.dmem1[i], inst_simd_top.inst_pe58_dmem.dmem0[i]
        };
       end

       $writememh("pe58.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe59_dmem.dmem3[i], inst_simd_top.inst_pe59_dmem.dmem2[i], inst_simd_top.inst_pe59_dmem.dmem1[i], inst_simd_top.inst_pe59_dmem.dmem0[i]
        };
       end

       $writememh("pe59.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe60_dmem.dmem3[i], inst_simd_top.inst_pe60_dmem.dmem2[i], inst_simd_top.inst_pe60_dmem.dmem1[i], inst_simd_top.inst_pe60_dmem.dmem0[i]
        };
       end

       $writememh("pe60.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe61_dmem.dmem3[i], inst_simd_top.inst_pe61_dmem.dmem2[i], inst_simd_top.inst_pe61_dmem.dmem1[i], inst_simd_top.inst_pe61_dmem.dmem0[i]
        };
       end

       $writememh("pe61.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe62_dmem.dmem3[i], inst_simd_top.inst_pe62_dmem.dmem2[i], inst_simd_top.inst_pe62_dmem.dmem1[i], inst_simd_top.inst_pe62_dmem.dmem0[i]
        };
       end

       $writememh("pe62.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe63_dmem.dmem3[i], inst_simd_top.inst_pe63_dmem.dmem2[i], inst_simd_top.inst_pe63_dmem.dmem1[i], inst_simd_top.inst_pe63_dmem.dmem0[i]
        };
       end

       $writememh("pe63.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe64_dmem.dmem3[i], inst_simd_top.inst_pe64_dmem.dmem2[i], inst_simd_top.inst_pe64_dmem.dmem1[i], inst_simd_top.inst_pe64_dmem.dmem0[i]
        };
       end

       $writememh("pe64.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe65_dmem.dmem3[i], inst_simd_top.inst_pe65_dmem.dmem2[i], inst_simd_top.inst_pe65_dmem.dmem1[i], inst_simd_top.inst_pe65_dmem.dmem0[i]
        };
       end

       $writememh("pe65.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe66_dmem.dmem3[i], inst_simd_top.inst_pe66_dmem.dmem2[i], inst_simd_top.inst_pe66_dmem.dmem1[i], inst_simd_top.inst_pe66_dmem.dmem0[i]
        };
       end

       $writememh("pe66.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe67_dmem.dmem3[i], inst_simd_top.inst_pe67_dmem.dmem2[i], inst_simd_top.inst_pe67_dmem.dmem1[i], inst_simd_top.inst_pe67_dmem.dmem0[i]
        };
       end

       $writememh("pe67.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe68_dmem.dmem3[i], inst_simd_top.inst_pe68_dmem.dmem2[i], inst_simd_top.inst_pe68_dmem.dmem1[i], inst_simd_top.inst_pe68_dmem.dmem0[i]
        };
       end

       $writememh("pe68.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe69_dmem.dmem3[i], inst_simd_top.inst_pe69_dmem.dmem2[i], inst_simd_top.inst_pe69_dmem.dmem1[i], inst_simd_top.inst_pe69_dmem.dmem0[i]
        };
       end

       $writememh("pe69.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe70_dmem.dmem3[i], inst_simd_top.inst_pe70_dmem.dmem2[i], inst_simd_top.inst_pe70_dmem.dmem1[i], inst_simd_top.inst_pe70_dmem.dmem0[i]
        };
       end

       $writememh("pe70.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe71_dmem.dmem3[i], inst_simd_top.inst_pe71_dmem.dmem2[i], inst_simd_top.inst_pe71_dmem.dmem1[i], inst_simd_top.inst_pe71_dmem.dmem0[i]
        };
       end

       $writememh("pe71.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe72_dmem.dmem3[i], inst_simd_top.inst_pe72_dmem.dmem2[i], inst_simd_top.inst_pe72_dmem.dmem1[i], inst_simd_top.inst_pe72_dmem.dmem0[i]
        };
       end

       $writememh("pe72.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe73_dmem.dmem3[i], inst_simd_top.inst_pe73_dmem.dmem2[i], inst_simd_top.inst_pe73_dmem.dmem1[i], inst_simd_top.inst_pe73_dmem.dmem0[i]
        };
       end

       $writememh("pe73.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe74_dmem.dmem3[i], inst_simd_top.inst_pe74_dmem.dmem2[i], inst_simd_top.inst_pe74_dmem.dmem1[i], inst_simd_top.inst_pe74_dmem.dmem0[i]
        };
       end

       $writememh("pe74.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe75_dmem.dmem3[i], inst_simd_top.inst_pe75_dmem.dmem2[i], inst_simd_top.inst_pe75_dmem.dmem1[i], inst_simd_top.inst_pe75_dmem.dmem0[i]
        };
       end

       $writememh("pe75.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe76_dmem.dmem3[i], inst_simd_top.inst_pe76_dmem.dmem2[i], inst_simd_top.inst_pe76_dmem.dmem1[i], inst_simd_top.inst_pe76_dmem.dmem0[i]
        };
       end

       $writememh("pe76.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe77_dmem.dmem3[i], inst_simd_top.inst_pe77_dmem.dmem2[i], inst_simd_top.inst_pe77_dmem.dmem1[i], inst_simd_top.inst_pe77_dmem.dmem0[i]
        };
       end

       $writememh("pe77.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe78_dmem.dmem3[i], inst_simd_top.inst_pe78_dmem.dmem2[i], inst_simd_top.inst_pe78_dmem.dmem1[i], inst_simd_top.inst_pe78_dmem.dmem0[i]
        };
       end

       $writememh("pe78.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe79_dmem.dmem3[i], inst_simd_top.inst_pe79_dmem.dmem2[i], inst_simd_top.inst_pe79_dmem.dmem1[i], inst_simd_top.inst_pe79_dmem.dmem0[i]
        };
       end

       $writememh("pe79.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe80_dmem.dmem3[i], inst_simd_top.inst_pe80_dmem.dmem2[i], inst_simd_top.inst_pe80_dmem.dmem1[i], inst_simd_top.inst_pe80_dmem.dmem0[i]
        };
       end

       $writememh("pe80.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe81_dmem.dmem3[i], inst_simd_top.inst_pe81_dmem.dmem2[i], inst_simd_top.inst_pe81_dmem.dmem1[i], inst_simd_top.inst_pe81_dmem.dmem0[i]
        };
       end

       $writememh("pe81.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe82_dmem.dmem3[i], inst_simd_top.inst_pe82_dmem.dmem2[i], inst_simd_top.inst_pe82_dmem.dmem1[i], inst_simd_top.inst_pe82_dmem.dmem0[i]
        };
       end

       $writememh("pe82.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe83_dmem.dmem3[i], inst_simd_top.inst_pe83_dmem.dmem2[i], inst_simd_top.inst_pe83_dmem.dmem1[i], inst_simd_top.inst_pe83_dmem.dmem0[i]
        };
       end

       $writememh("pe83.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe84_dmem.dmem3[i], inst_simd_top.inst_pe84_dmem.dmem2[i], inst_simd_top.inst_pe84_dmem.dmem1[i], inst_simd_top.inst_pe84_dmem.dmem0[i]
        };
       end

       $writememh("pe84.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe85_dmem.dmem3[i], inst_simd_top.inst_pe85_dmem.dmem2[i], inst_simd_top.inst_pe85_dmem.dmem1[i], inst_simd_top.inst_pe85_dmem.dmem0[i]
        };
       end

       $writememh("pe85.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe86_dmem.dmem3[i], inst_simd_top.inst_pe86_dmem.dmem2[i], inst_simd_top.inst_pe86_dmem.dmem1[i], inst_simd_top.inst_pe86_dmem.dmem0[i]
        };
       end

       $writememh("pe86.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe87_dmem.dmem3[i], inst_simd_top.inst_pe87_dmem.dmem2[i], inst_simd_top.inst_pe87_dmem.dmem1[i], inst_simd_top.inst_pe87_dmem.dmem0[i]
        };
       end

       $writememh("pe87.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe88_dmem.dmem3[i], inst_simd_top.inst_pe88_dmem.dmem2[i], inst_simd_top.inst_pe88_dmem.dmem1[i], inst_simd_top.inst_pe88_dmem.dmem0[i]
        };
       end

       $writememh("pe88.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe89_dmem.dmem3[i], inst_simd_top.inst_pe89_dmem.dmem2[i], inst_simd_top.inst_pe89_dmem.dmem1[i], inst_simd_top.inst_pe89_dmem.dmem0[i]
        };
       end

       $writememh("pe89.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe90_dmem.dmem3[i], inst_simd_top.inst_pe90_dmem.dmem2[i], inst_simd_top.inst_pe90_dmem.dmem1[i], inst_simd_top.inst_pe90_dmem.dmem0[i]
        };
       end

       $writememh("pe90.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe91_dmem.dmem3[i], inst_simd_top.inst_pe91_dmem.dmem2[i], inst_simd_top.inst_pe91_dmem.dmem1[i], inst_simd_top.inst_pe91_dmem.dmem0[i]
        };
       end

       $writememh("pe91.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe92_dmem.dmem3[i], inst_simd_top.inst_pe92_dmem.dmem2[i], inst_simd_top.inst_pe92_dmem.dmem1[i], inst_simd_top.inst_pe92_dmem.dmem0[i]
        };
       end

       $writememh("pe92.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe93_dmem.dmem3[i], inst_simd_top.inst_pe93_dmem.dmem2[i], inst_simd_top.inst_pe93_dmem.dmem1[i], inst_simd_top.inst_pe93_dmem.dmem0[i]
        };
       end

       $writememh("pe93.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe94_dmem.dmem3[i], inst_simd_top.inst_pe94_dmem.dmem2[i], inst_simd_top.inst_pe94_dmem.dmem1[i], inst_simd_top.inst_pe94_dmem.dmem0[i]
        };
       end

       $writememh("pe94.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe95_dmem.dmem3[i], inst_simd_top.inst_pe95_dmem.dmem2[i], inst_simd_top.inst_pe95_dmem.dmem1[i], inst_simd_top.inst_pe95_dmem.dmem0[i]
        };
       end

       $writememh("pe95.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe96_dmem.dmem3[i], inst_simd_top.inst_pe96_dmem.dmem2[i], inst_simd_top.inst_pe96_dmem.dmem1[i], inst_simd_top.inst_pe96_dmem.dmem0[i]
        };
       end

       $writememh("pe96.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe97_dmem.dmem3[i], inst_simd_top.inst_pe97_dmem.dmem2[i], inst_simd_top.inst_pe97_dmem.dmem1[i], inst_simd_top.inst_pe97_dmem.dmem0[i]
        };
       end

       $writememh("pe97.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe98_dmem.dmem3[i], inst_simd_top.inst_pe98_dmem.dmem2[i], inst_simd_top.inst_pe98_dmem.dmem1[i], inst_simd_top.inst_pe98_dmem.dmem0[i]
        };
       end

       $writememh("pe98.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe99_dmem.dmem3[i], inst_simd_top.inst_pe99_dmem.dmem2[i], inst_simd_top.inst_pe99_dmem.dmem1[i], inst_simd_top.inst_pe99_dmem.dmem0[i]
        };
       end

       $writememh("pe99.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe100_dmem.dmem3[i], inst_simd_top.inst_pe100_dmem.dmem2[i], inst_simd_top.inst_pe100_dmem.dmem1[i], inst_simd_top.inst_pe100_dmem.dmem0[i]
        };
       end

       $writememh("pe100.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe101_dmem.dmem3[i], inst_simd_top.inst_pe101_dmem.dmem2[i], inst_simd_top.inst_pe101_dmem.dmem1[i], inst_simd_top.inst_pe101_dmem.dmem0[i]
        };
       end

       $writememh("pe101.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe102_dmem.dmem3[i], inst_simd_top.inst_pe102_dmem.dmem2[i], inst_simd_top.inst_pe102_dmem.dmem1[i], inst_simd_top.inst_pe102_dmem.dmem0[i]
        };
       end

       $writememh("pe102.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe103_dmem.dmem3[i], inst_simd_top.inst_pe103_dmem.dmem2[i], inst_simd_top.inst_pe103_dmem.dmem1[i], inst_simd_top.inst_pe103_dmem.dmem0[i]
        };
       end

       $writememh("pe103.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe104_dmem.dmem3[i], inst_simd_top.inst_pe104_dmem.dmem2[i], inst_simd_top.inst_pe104_dmem.dmem1[i], inst_simd_top.inst_pe104_dmem.dmem0[i]
        };
       end

       $writememh("pe104.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe105_dmem.dmem3[i], inst_simd_top.inst_pe105_dmem.dmem2[i], inst_simd_top.inst_pe105_dmem.dmem1[i], inst_simd_top.inst_pe105_dmem.dmem0[i]
        };
       end

       $writememh("pe105.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe106_dmem.dmem3[i], inst_simd_top.inst_pe106_dmem.dmem2[i], inst_simd_top.inst_pe106_dmem.dmem1[i], inst_simd_top.inst_pe106_dmem.dmem0[i]
        };
       end

       $writememh("pe106.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe107_dmem.dmem3[i], inst_simd_top.inst_pe107_dmem.dmem2[i], inst_simd_top.inst_pe107_dmem.dmem1[i], inst_simd_top.inst_pe107_dmem.dmem0[i]
        };
       end

       $writememh("pe107.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe108_dmem.dmem3[i], inst_simd_top.inst_pe108_dmem.dmem2[i], inst_simd_top.inst_pe108_dmem.dmem1[i], inst_simd_top.inst_pe108_dmem.dmem0[i]
        };
       end

       $writememh("pe108.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe109_dmem.dmem3[i], inst_simd_top.inst_pe109_dmem.dmem2[i], inst_simd_top.inst_pe109_dmem.dmem1[i], inst_simd_top.inst_pe109_dmem.dmem0[i]
        };
       end

       $writememh("pe109.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe110_dmem.dmem3[i], inst_simd_top.inst_pe110_dmem.dmem2[i], inst_simd_top.inst_pe110_dmem.dmem1[i], inst_simd_top.inst_pe110_dmem.dmem0[i]
        };
       end

       $writememh("pe110.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe111_dmem.dmem3[i], inst_simd_top.inst_pe111_dmem.dmem2[i], inst_simd_top.inst_pe111_dmem.dmem1[i], inst_simd_top.inst_pe111_dmem.dmem0[i]
        };
       end

       $writememh("pe111.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe112_dmem.dmem3[i], inst_simd_top.inst_pe112_dmem.dmem2[i], inst_simd_top.inst_pe112_dmem.dmem1[i], inst_simd_top.inst_pe112_dmem.dmem0[i]
        };
       end

       $writememh("pe112.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe113_dmem.dmem3[i], inst_simd_top.inst_pe113_dmem.dmem2[i], inst_simd_top.inst_pe113_dmem.dmem1[i], inst_simd_top.inst_pe113_dmem.dmem0[i]
        };
       end

       $writememh("pe113.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe114_dmem.dmem3[i], inst_simd_top.inst_pe114_dmem.dmem2[i], inst_simd_top.inst_pe114_dmem.dmem1[i], inst_simd_top.inst_pe114_dmem.dmem0[i]
        };
       end

       $writememh("pe114.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe115_dmem.dmem3[i], inst_simd_top.inst_pe115_dmem.dmem2[i], inst_simd_top.inst_pe115_dmem.dmem1[i], inst_simd_top.inst_pe115_dmem.dmem0[i]
        };
       end

       $writememh("pe115.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe116_dmem.dmem3[i], inst_simd_top.inst_pe116_dmem.dmem2[i], inst_simd_top.inst_pe116_dmem.dmem1[i], inst_simd_top.inst_pe116_dmem.dmem0[i]
        };
       end

       $writememh("pe116.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe117_dmem.dmem3[i], inst_simd_top.inst_pe117_dmem.dmem2[i], inst_simd_top.inst_pe117_dmem.dmem1[i], inst_simd_top.inst_pe117_dmem.dmem0[i]
        };
       end

       $writememh("pe117.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe118_dmem.dmem3[i], inst_simd_top.inst_pe118_dmem.dmem2[i], inst_simd_top.inst_pe118_dmem.dmem1[i], inst_simd_top.inst_pe118_dmem.dmem0[i]
        };
       end

       $writememh("pe118.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe119_dmem.dmem3[i], inst_simd_top.inst_pe119_dmem.dmem2[i], inst_simd_top.inst_pe119_dmem.dmem1[i], inst_simd_top.inst_pe119_dmem.dmem0[i]
        };
       end

       $writememh("pe119.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe120_dmem.dmem3[i], inst_simd_top.inst_pe120_dmem.dmem2[i], inst_simd_top.inst_pe120_dmem.dmem1[i], inst_simd_top.inst_pe120_dmem.dmem0[i]
        };
       end

       $writememh("pe120.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe121_dmem.dmem3[i], inst_simd_top.inst_pe121_dmem.dmem2[i], inst_simd_top.inst_pe121_dmem.dmem1[i], inst_simd_top.inst_pe121_dmem.dmem0[i]
        };
       end

       $writememh("pe121.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe122_dmem.dmem3[i], inst_simd_top.inst_pe122_dmem.dmem2[i], inst_simd_top.inst_pe122_dmem.dmem1[i], inst_simd_top.inst_pe122_dmem.dmem0[i]
        };
       end

       $writememh("pe122.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe123_dmem.dmem3[i], inst_simd_top.inst_pe123_dmem.dmem2[i], inst_simd_top.inst_pe123_dmem.dmem1[i], inst_simd_top.inst_pe123_dmem.dmem0[i]
        };
       end

       $writememh("pe123.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe124_dmem.dmem3[i], inst_simd_top.inst_pe124_dmem.dmem2[i], inst_simd_top.inst_pe124_dmem.dmem1[i], inst_simd_top.inst_pe124_dmem.dmem0[i]
        };
       end

       $writememh("pe124.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe125_dmem.dmem3[i], inst_simd_top.inst_pe125_dmem.dmem2[i], inst_simd_top.inst_pe125_dmem.dmem1[i], inst_simd_top.inst_pe125_dmem.dmem0[i]
        };
       end

       $writememh("pe125.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe126_dmem.dmem3[i], inst_simd_top.inst_pe126_dmem.dmem2[i], inst_simd_top.inst_pe126_dmem.dmem1[i], inst_simd_top.inst_pe126_dmem.dmem0[i]
        };
       end

       $writememh("pe126.dmem.dump", PE_DMEM_tmp);

       for (i=0; i<`DEF_PE_DMEM_SIZE; i=i+1) begin
        PE_DMEM_tmp[i] = {inst_simd_top.inst_pe127_dmem.dmem3[i], inst_simd_top.inst_pe127_dmem.dmem2[i], inst_simd_top.inst_pe127_dmem.dmem1[i], inst_simd_top.inst_pe127_dmem.dmem0[i]
        };
       end

       $writememh("pe127.dmem.dump", PE_DMEM_tmp);

       
       $finish;
     end
  // end of initial

  // core reset: active high
  assign wCore_Reset = ~( rReset && rIMEM_Configure_Done && rCP_DMEM_Configure_Done && rPE_DMEM_Configure_Done );

  simd_top inst_simd_top (
    .iClk                          ( rClk                      ), // system clock, positive-edge trigger
    .iReset                        ( wCore_Reset               ), // global synchronous reset signal, Active high

    .oIF_ID_PC                     ( wPC                       ), // current PC for debug
    .oTask_Finished                ( wTask_Finished            ), // indicate the end of the program

    // Instruction Memory
    .iBus_CP_IMEM_Valid            ( rBus_IMEM_Valid           ), // cp ins. memory access valid
    .iBus_CP_IMEM_Address          ( rBus_IMEM_Address         ), // cp ins. memory access address
    .iBus_CP_IMEM_Write_Data       ( rBus_IMEM_Write_Data[(`DEF_CP_INS_WIDTH+3):0] ), // cp ins. memory write data
    .iBus_CP_IMEM_Write_Enable     ( rBus_IMEM_Write_Enable    ), // cp ins. memory write enable
    .oBus_CP_IMEM_Read_Data        ( wBus_CP_IMEM_Read_Data    ), // cp ins. memory read data

    .iBus_PE_IMEM_Valid            ( rBus_IMEM_Valid           ), // pe ins. memory access valid
    .iBus_PE_IMEM_Address          ( rBus_IMEM_Address         ), // pe ins. memory access address
    .iBus_PE_IMEM_Write_Data       ( rBus_IMEM_Write_Data[(`DEF_PE_INS_WIDTH+4)+32:32] ), // pe ins. memory write data
    .iBus_PE_IMEM_Write_Enable     ( rBus_IMEM_Write_Enable    ), // pe ins. memory write enable
    .oBus_PE_IMEM_Read_Data        ( wBus_PE_IMEM_Read_Data    ), // pe ins. memory read data

    // Data Memory
    .iBus_CP_DMEM_Valid            ( rBus_CP_DMEM_Valid        ), // cp data memory access valid
    .iBus_CP_DMEM_Address          ( {rBus_CP_DMEM_Address, 2'b0} ), // cp data memory access address
    .iBus_CP_DMEM_Write_Data       ( rBus_CP_DMEM_Write_Data   ), // cp data memory write data
    .iBus_CP_DMEM_Write_Enable     ( rBus_CP_DMEM_Write_Enable ), // cp data memory write enable
    .oBus_CP_DMEM_Read_Data        ( wBus_CP_DMEM_Read_Data    ), // cp data memory read data

    .iBus_PE_DMEM_Valid            ( {`DEF_PE_NUM{rBus_PE_DMEM_Valid}} ), // pe data memory access valid
    .iBus_PE_DMEM_Address          ( {`DEF_PE_NUM{rBus_PE_DMEM_Address, 2'b0}} ), // pe data memory access address
    .iBus_PE_DMEM_Write_Data       ( rBus_PE_DMEM_Write_Data  ), // pe data memory write data
    .iBus_PE_DMEM_Write_Enable     ( {`DEF_PE_NUM{rBus_PE_DMEM_Write_Enable}} ), // pe data memory write enable
    .oBus_PE_DMEM_Read_Data        ( wBus_PE_DMEM_Read_Data   )  // pe data memory read data
  );


endmodule