library verilog;
use verilog.vl_types.all;
entity simd_top_testbench is
end simd_top_testbench;
