library verilog;
use verilog.vl_types.all;
entity core_top is
    port(
        iClk            : in     vl_logic;
        iReset          : in     vl_logic;
        oIF_ID_PC       : out    vl_logic_vector(16 downto 0);
        oTask_Finished  : out    vl_logic;
        oIF_IMEM_Address: out    vl_logic_vector(16 downto 0);
        iIMEM_CP_Instruction: in     vl_logic_vector(27 downto 0);
        oCP_DMEM_Valid  : out    vl_logic;
        oCP_AGU_DMEM_Write_Enable: out    vl_logic;
        oCP_AGU_DMEM_Read_Enable: out    vl_logic;
        oCP_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oCP_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oCP_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iCP_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE0_DMEM_Valid : out    vl_logic;
        oPE0_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE0_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE0_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE0_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE0_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE0_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE1_DMEM_Valid : out    vl_logic;
        oPE1_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE1_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE1_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE1_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE1_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE1_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE2_DMEM_Valid : out    vl_logic;
        oPE2_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE2_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE2_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE2_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE2_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE2_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE3_DMEM_Valid : out    vl_logic;
        oPE3_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE3_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE3_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE3_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE3_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE3_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE4_DMEM_Valid : out    vl_logic;
        oPE4_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE4_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE4_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE4_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE4_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE4_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE5_DMEM_Valid : out    vl_logic;
        oPE5_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE5_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE5_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE5_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE5_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE5_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE6_DMEM_Valid : out    vl_logic;
        oPE6_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE6_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE6_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE6_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE6_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE6_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE7_DMEM_Valid : out    vl_logic;
        oPE7_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE7_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE7_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE7_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE7_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE7_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE8_DMEM_Valid : out    vl_logic;
        oPE8_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE8_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE8_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE8_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE8_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE8_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE9_DMEM_Valid : out    vl_logic;
        oPE9_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE9_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE9_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE9_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE9_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE9_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE10_DMEM_Valid: out    vl_logic;
        oPE10_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE10_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE10_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE10_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE10_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE10_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE11_DMEM_Valid: out    vl_logic;
        oPE11_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE11_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE11_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE11_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE11_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE11_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE12_DMEM_Valid: out    vl_logic;
        oPE12_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE12_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE12_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE12_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE12_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE12_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE13_DMEM_Valid: out    vl_logic;
        oPE13_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE13_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE13_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE13_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE13_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE13_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE14_DMEM_Valid: out    vl_logic;
        oPE14_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE14_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE14_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE14_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE14_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE14_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE15_DMEM_Valid: out    vl_logic;
        oPE15_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE15_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE15_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE15_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE15_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE15_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE16_DMEM_Valid: out    vl_logic;
        oPE16_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE16_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE16_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE16_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE16_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE16_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE17_DMEM_Valid: out    vl_logic;
        oPE17_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE17_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE17_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE17_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE17_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE17_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE18_DMEM_Valid: out    vl_logic;
        oPE18_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE18_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE18_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE18_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE18_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE18_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE19_DMEM_Valid: out    vl_logic;
        oPE19_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE19_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE19_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE19_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE19_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE19_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE20_DMEM_Valid: out    vl_logic;
        oPE20_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE20_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE20_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE20_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE20_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE20_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE21_DMEM_Valid: out    vl_logic;
        oPE21_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE21_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE21_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE21_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE21_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE21_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE22_DMEM_Valid: out    vl_logic;
        oPE22_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE22_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE22_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE22_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE22_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE22_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE23_DMEM_Valid: out    vl_logic;
        oPE23_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE23_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE23_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE23_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE23_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE23_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE24_DMEM_Valid: out    vl_logic;
        oPE24_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE24_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE24_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE24_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE24_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE24_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE25_DMEM_Valid: out    vl_logic;
        oPE25_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE25_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE25_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE25_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE25_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE25_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE26_DMEM_Valid: out    vl_logic;
        oPE26_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE26_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE26_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE26_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE26_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE26_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE27_DMEM_Valid: out    vl_logic;
        oPE27_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE27_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE27_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE27_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE27_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE27_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE28_DMEM_Valid: out    vl_logic;
        oPE28_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE28_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE28_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE28_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE28_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE28_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE29_DMEM_Valid: out    vl_logic;
        oPE29_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE29_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE29_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE29_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE29_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE29_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE30_DMEM_Valid: out    vl_logic;
        oPE30_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE30_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE30_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE30_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE30_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE30_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE31_DMEM_Valid: out    vl_logic;
        oPE31_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE31_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE31_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE31_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE31_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE31_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE32_DMEM_Valid: out    vl_logic;
        oPE32_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE32_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE32_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE32_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE32_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE32_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE33_DMEM_Valid: out    vl_logic;
        oPE33_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE33_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE33_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE33_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE33_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE33_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE34_DMEM_Valid: out    vl_logic;
        oPE34_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE34_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE34_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE34_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE34_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE34_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE35_DMEM_Valid: out    vl_logic;
        oPE35_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE35_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE35_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE35_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE35_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE35_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE36_DMEM_Valid: out    vl_logic;
        oPE36_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE36_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE36_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE36_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE36_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE36_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE37_DMEM_Valid: out    vl_logic;
        oPE37_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE37_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE37_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE37_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE37_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE37_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE38_DMEM_Valid: out    vl_logic;
        oPE38_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE38_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE38_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE38_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE38_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE38_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE39_DMEM_Valid: out    vl_logic;
        oPE39_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE39_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE39_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE39_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE39_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE39_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE40_DMEM_Valid: out    vl_logic;
        oPE40_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE40_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE40_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE40_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE40_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE40_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE41_DMEM_Valid: out    vl_logic;
        oPE41_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE41_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE41_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE41_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE41_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE41_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE42_DMEM_Valid: out    vl_logic;
        oPE42_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE42_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE42_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE42_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE42_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE42_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE43_DMEM_Valid: out    vl_logic;
        oPE43_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE43_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE43_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE43_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE43_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE43_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE44_DMEM_Valid: out    vl_logic;
        oPE44_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE44_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE44_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE44_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE44_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE44_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE45_DMEM_Valid: out    vl_logic;
        oPE45_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE45_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE45_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE45_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE45_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE45_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE46_DMEM_Valid: out    vl_logic;
        oPE46_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE46_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE46_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE46_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE46_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE46_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE47_DMEM_Valid: out    vl_logic;
        oPE47_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE47_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE47_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE47_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE47_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE47_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE48_DMEM_Valid: out    vl_logic;
        oPE48_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE48_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE48_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE48_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE48_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE48_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE49_DMEM_Valid: out    vl_logic;
        oPE49_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE49_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE49_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE49_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE49_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE49_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE50_DMEM_Valid: out    vl_logic;
        oPE50_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE50_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE50_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE50_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE50_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE50_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE51_DMEM_Valid: out    vl_logic;
        oPE51_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE51_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE51_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE51_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE51_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE51_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE52_DMEM_Valid: out    vl_logic;
        oPE52_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE52_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE52_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE52_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE52_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE52_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE53_DMEM_Valid: out    vl_logic;
        oPE53_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE53_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE53_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE53_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE53_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE53_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE54_DMEM_Valid: out    vl_logic;
        oPE54_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE54_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE54_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE54_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE54_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE54_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE55_DMEM_Valid: out    vl_logic;
        oPE55_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE55_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE55_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE55_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE55_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE55_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE56_DMEM_Valid: out    vl_logic;
        oPE56_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE56_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE56_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE56_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE56_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE56_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE57_DMEM_Valid: out    vl_logic;
        oPE57_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE57_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE57_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE57_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE57_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE57_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE58_DMEM_Valid: out    vl_logic;
        oPE58_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE58_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE58_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE58_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE58_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE58_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE59_DMEM_Valid: out    vl_logic;
        oPE59_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE59_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE59_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE59_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE59_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE59_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE60_DMEM_Valid: out    vl_logic;
        oPE60_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE60_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE60_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE60_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE60_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE60_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE61_DMEM_Valid: out    vl_logic;
        oPE61_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE61_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE61_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE61_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE61_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE61_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE62_DMEM_Valid: out    vl_logic;
        oPE62_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE62_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE62_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE62_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE62_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE62_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE63_DMEM_Valid: out    vl_logic;
        oPE63_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE63_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE63_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE63_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE63_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE63_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE64_DMEM_Valid: out    vl_logic;
        oPE64_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE64_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE64_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE64_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE64_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE64_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE65_DMEM_Valid: out    vl_logic;
        oPE65_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE65_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE65_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE65_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE65_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE65_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE66_DMEM_Valid: out    vl_logic;
        oPE66_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE66_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE66_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE66_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE66_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE66_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE67_DMEM_Valid: out    vl_logic;
        oPE67_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE67_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE67_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE67_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE67_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE67_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE68_DMEM_Valid: out    vl_logic;
        oPE68_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE68_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE68_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE68_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE68_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE68_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE69_DMEM_Valid: out    vl_logic;
        oPE69_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE69_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE69_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE69_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE69_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE69_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE70_DMEM_Valid: out    vl_logic;
        oPE70_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE70_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE70_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE70_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE70_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE70_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE71_DMEM_Valid: out    vl_logic;
        oPE71_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE71_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE71_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE71_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE71_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE71_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE72_DMEM_Valid: out    vl_logic;
        oPE72_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE72_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE72_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE72_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE72_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE72_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE73_DMEM_Valid: out    vl_logic;
        oPE73_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE73_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE73_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE73_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE73_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE73_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE74_DMEM_Valid: out    vl_logic;
        oPE74_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE74_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE74_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE74_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE74_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE74_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE75_DMEM_Valid: out    vl_logic;
        oPE75_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE75_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE75_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE75_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE75_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE75_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE76_DMEM_Valid: out    vl_logic;
        oPE76_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE76_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE76_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE76_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE76_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE76_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE77_DMEM_Valid: out    vl_logic;
        oPE77_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE77_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE77_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE77_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE77_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE77_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE78_DMEM_Valid: out    vl_logic;
        oPE78_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE78_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE78_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE78_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE78_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE78_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE79_DMEM_Valid: out    vl_logic;
        oPE79_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE79_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE79_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE79_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE79_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE79_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE80_DMEM_Valid: out    vl_logic;
        oPE80_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE80_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE80_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE80_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE80_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE80_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE81_DMEM_Valid: out    vl_logic;
        oPE81_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE81_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE81_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE81_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE81_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE81_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE82_DMEM_Valid: out    vl_logic;
        oPE82_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE82_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE82_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE82_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE82_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE82_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE83_DMEM_Valid: out    vl_logic;
        oPE83_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE83_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE83_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE83_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE83_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE83_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE84_DMEM_Valid: out    vl_logic;
        oPE84_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE84_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE84_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE84_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE84_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE84_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE85_DMEM_Valid: out    vl_logic;
        oPE85_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE85_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE85_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE85_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE85_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE85_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE86_DMEM_Valid: out    vl_logic;
        oPE86_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE86_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE86_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE86_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE86_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE86_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE87_DMEM_Valid: out    vl_logic;
        oPE87_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE87_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE87_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE87_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE87_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE87_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE88_DMEM_Valid: out    vl_logic;
        oPE88_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE88_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE88_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE88_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE88_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE88_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE89_DMEM_Valid: out    vl_logic;
        oPE89_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE89_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE89_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE89_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE89_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE89_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE90_DMEM_Valid: out    vl_logic;
        oPE90_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE90_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE90_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE90_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE90_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE90_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE91_DMEM_Valid: out    vl_logic;
        oPE91_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE91_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE91_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE91_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE91_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE91_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE92_DMEM_Valid: out    vl_logic;
        oPE92_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE92_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE92_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE92_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE92_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE92_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE93_DMEM_Valid: out    vl_logic;
        oPE93_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE93_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE93_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE93_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE93_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE93_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE94_DMEM_Valid: out    vl_logic;
        oPE94_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE94_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE94_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE94_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE94_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE94_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE95_DMEM_Valid: out    vl_logic;
        oPE95_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE95_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE95_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE95_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE95_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE95_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE96_DMEM_Valid: out    vl_logic;
        oPE96_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE96_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE96_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE96_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE96_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE96_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE97_DMEM_Valid: out    vl_logic;
        oPE97_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE97_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE97_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE97_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE97_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE97_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE98_DMEM_Valid: out    vl_logic;
        oPE98_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE98_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE98_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE98_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE98_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE98_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE99_DMEM_Valid: out    vl_logic;
        oPE99_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE99_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE99_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE99_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE99_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE99_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE100_DMEM_Valid: out    vl_logic;
        oPE100_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE100_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE100_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE100_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE100_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE100_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE101_DMEM_Valid: out    vl_logic;
        oPE101_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE101_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE101_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE101_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE101_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE101_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE102_DMEM_Valid: out    vl_logic;
        oPE102_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE102_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE102_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE102_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE102_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE102_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE103_DMEM_Valid: out    vl_logic;
        oPE103_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE103_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE103_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE103_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE103_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE103_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE104_DMEM_Valid: out    vl_logic;
        oPE104_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE104_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE104_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE104_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE104_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE104_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE105_DMEM_Valid: out    vl_logic;
        oPE105_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE105_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE105_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE105_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE105_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE105_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE106_DMEM_Valid: out    vl_logic;
        oPE106_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE106_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE106_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE106_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE106_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE106_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE107_DMEM_Valid: out    vl_logic;
        oPE107_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE107_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE107_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE107_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE107_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE107_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE108_DMEM_Valid: out    vl_logic;
        oPE108_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE108_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE108_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE108_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE108_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE108_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE109_DMEM_Valid: out    vl_logic;
        oPE109_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE109_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE109_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE109_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE109_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE109_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE110_DMEM_Valid: out    vl_logic;
        oPE110_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE110_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE110_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE110_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE110_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE110_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE111_DMEM_Valid: out    vl_logic;
        oPE111_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE111_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE111_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE111_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE111_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE111_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE112_DMEM_Valid: out    vl_logic;
        oPE112_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE112_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE112_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE112_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE112_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE112_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE113_DMEM_Valid: out    vl_logic;
        oPE113_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE113_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE113_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE113_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE113_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE113_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE114_DMEM_Valid: out    vl_logic;
        oPE114_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE114_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE114_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE114_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE114_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE114_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE115_DMEM_Valid: out    vl_logic;
        oPE115_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE115_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE115_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE115_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE115_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE115_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE116_DMEM_Valid: out    vl_logic;
        oPE116_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE116_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE116_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE116_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE116_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE116_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE117_DMEM_Valid: out    vl_logic;
        oPE117_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE117_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE117_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE117_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE117_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE117_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE118_DMEM_Valid: out    vl_logic;
        oPE118_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE118_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE118_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE118_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE118_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE118_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE119_DMEM_Valid: out    vl_logic;
        oPE119_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE119_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE119_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE119_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE119_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE119_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE120_DMEM_Valid: out    vl_logic;
        oPE120_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE120_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE120_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE120_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE120_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE120_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE121_DMEM_Valid: out    vl_logic;
        oPE121_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE121_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE121_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE121_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE121_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE121_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE122_DMEM_Valid: out    vl_logic;
        oPE122_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE122_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE122_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE122_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE122_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE122_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE123_DMEM_Valid: out    vl_logic;
        oPE123_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE123_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE123_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE123_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE123_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE123_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE124_DMEM_Valid: out    vl_logic;
        oPE124_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE124_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE124_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE124_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE124_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE124_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE125_DMEM_Valid: out    vl_logic;
        oPE125_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE125_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE125_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE125_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE125_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE125_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE126_DMEM_Valid: out    vl_logic;
        oPE126_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE126_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE126_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE126_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE126_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE126_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        oPE127_DMEM_Valid: out    vl_logic;
        oPE127_AGU_DMEM_Write_Enable: out    vl_logic;
        oPE127_AGU_DMEM_Read_Enable: out    vl_logic;
        oPE127_AGU_DMEM_Byte_Select: out    vl_logic_vector(3 downto 0);
        oPE127_AGU_DMEM_Address: out    vl_logic_vector(10 downto 0);
        oPE127_AGU_DMEM_Write_Data: out    vl_logic_vector(31 downto 0);
        iPE127_DMEM_EX_Data: in     vl_logic_vector(31 downto 0);
        iIMEM_PE_Instruction: in     vl_logic_vector(28 downto 0)
    );
end core_top;
